module truncator (
input [127:0]a,
output reg [51:0]b,
output reg setzero
);
//assign setzero = 0;
always@(a)
begin
	if(a[127]) b[51:0] = a[127:76];
	else if(a[126]) b[51:0] = a[126:75];
	else if(a[125]) b[51:0] = a[125:74];
	else if(a[124]) b[51:0] = a[124:73];

	else if(a[123]) b[51:0] = a[123:72];
	else if(a[122]) b[51:0] = a[122:71];
	else if(a[121]) b[51:0] = a[121:70];
	else if(a[120]) b[51:0] = a[120:69];
	else if(a[119]) b[51:0] = a[119:68];
	else if(a[118]) b[51:0] = a[118:67];
	else if(a[117]) b[51:0] = a[117:66];
	else if(a[116]) b[51:0] = a[116:65];
	else if(a[115]) b[51:0] = a[115:64];
	else if(a[114]) b[51:0] = a[114:63];
	else if(a[113]) b[51:0] = a[113:62];
	else if(a[112]) b[51:0] = a[112:61];
	else if(a[111]) b[51:0] = a[111:60];
	else if(a[110]) b[51:0] = a[110:59];
	else if(a[109]) b[51:0] = a[109:58];
	else if(a[108]) b[51:0] = a[108:57];
	else if(a[107]) b[51:0] = a[107:56];
	else if(a[106]) b[51:0] = a[106:55];
	else if(a[105]) b[51:0] = a[105:54];
	else if(a[104]) b[51:0] = a[104:53];
	else if(a[103]) b[51:0] = a[103:52];
	else if(a[102]) b[51:0] = a[102:51];
	else if(a[101]) b[51:0] = a[101:50];
	else if(a[100]) b[51:0] = a[100:49];


	else if(a[99]) b[51:0] = a[99:48];
	else if(a[98]) b[51:0] = a[98:47];
	else if(a[97]) b[51:0] = a[97:46];
	else if(a[96]) b[51:0] = a[96:45];
	else if(a[95]) b[51:0] = a[95:44];
	else if(a[94]) b[51:0] = a[94:43];
	else if(a[93]) b[51:0] = a[93:42];
	else if(a[92]) b[51:0] = a[92:41];
	else if(a[91]) b[51:0] = a[91:40];
	else if(a[90]) b[51:0] = a[90:39];
	
	else if(a[89]) b[51:0] = a[89:38];
	else if(a[88]) b[51:0] = a[88:37];
	else if(a[87]) b[51:0] = a[87:36];
	else if(a[86]) b[51:0] = a[86:35];
	else if(a[85]) b[51:0] = a[85:34];
	else if(a[84]) b[51:0] = a[84:33];
	else if(a[83]) b[51:0] = a[83:32];
	else if(a[82]) b[51:0] = a[82:31];
	else if(a[81]) b[51:0] = a[81:30];
	else if(a[80]) b[51:0] = a[80:29];

	else if(a[79]) b[51:0] = a[79:28];
	else if(a[78]) b[51:0] = a[78:27];
	else if(a[77]) b[51:0] = a[77:26];
	else if(a[76]) b[51:0] = a[76:25];
	else if(a[75]) b[51:0] = a[75:24];
	else if(a[74]) b[51:0] = a[74:23];
	else if(a[73]) b[51:0] = a[73:22];
	else if(a[72]) b[51:0] = a[72:21];
	else if(a[71]) b[51:0] = a[71:20];
	else if(a[70]) b[51:0] = a[70:19];
	
	else if(a[69]) b[51:0] = a[69:18];
	else if(a[68]) b[51:0] = a[68:17];
	else if(a[67]) b[51:0] = a[67:16];
	else if(a[66]) b[51:0] = a[66:15];
	else if(a[65]) b[51:0] = a[65:14];
	else if(a[64]) b[51:0] = a[64:13];
	else if(a[63]) b[51:0] = a[63:12];
	else if(a[62]) b[51:0] = a[62:11];
	else if(a[61]) b[51:0] = a[61:10];
	else if(a[60]) b[51:0] = a[60:9];
	
	else if(a[59]) b[51:0] = a[59:8];
	else if(a[58]) b[51:0] = a[58:7];
	else if(a[57]) b[51:0] = a[57:6];
	else if(a[56]) b[51:0] = a[56:5];
	else if(a[55]) b[51:0] = a[55:4];
	else if(a[54]) b[51:0] = a[54:3];
	else if(a[53]) b[51:0] = a[53:2];
	else if(a[52]) b[51:0] = a[52:1];
	else if(a[51]) b[51:0] = a[51:0];
	else if(a[50]) b[51:0] = {a[50:0],1'b0};
	
	
	else if(a[49]) b[51:0] = {a[49:0],2'b0};
	else if(a[48]) b[51:0] = {a[48:0],3'b0};
	else if(a[47]) b[51:0] = {a[47:0],4'b0};
	else if(a[46]) b[51:0] = {a[46:0],5'b0};
	else if(a[45]) b[51:0] = {a[45:0],6'b0};
	else if(a[44]) b[51:0] = {a[44:0],7'b0};
	else if(a[43]) b[51:0] = {a[43:0],8'b0};
	else if(a[42]) b[51:0] = {a[42:0],9'b0};
	else if(a[41]) b[51:0] = {a[41:0],10'b0};
	else if(a[40]) b[51:0] = {a[40:0],11'b0};
	
	else if(a[39]) b[51:0] = {a[39:0],12'b0};
	else if(a[38]) b[51:0] = {a[38:0],13'b0};
	else if(a[37]) b[51:0] = {a[37:0],14'b0};
	else if(a[36]) b[51:0] = {a[36:0],15'b0};
	else if(a[35]) b[51:0] = {a[35:0],16'b0};
	else if(a[34]) b[51:0] = {a[34:0],17'b0};
	else if(a[33]) b[51:0] = {a[33:0],18'b0};
	else if(a[32]) b[51:0] = {a[32:0],19'b0};
	else if(a[31]) b[51:0] = {a[31:0],20'b0};
	else if(a[30]) b[51:0] = {a[30:0],21'b0};




	
	
	
	
	else if(a[29]) b[51:0] = {a[29:0],22'b0};
	else if(a[28]) b[51:0] = {a[28:0],23'b0};
	else if(a[27]) b[51:0] = {a[27:0],24'b0};
	else if(a[26]) b[51:0] = {a[26:0],25'b0};
	else if(a[25]) b[51:0] = {a[25:0],26'b0};
	else if(a[24]) b[51:0] = {a[24:0],27'b0};
	else if(a[23]) b[51:0] = {a[23:0],28'b0};
	else if(a[22]) b[51:0] = {a[22:0],29'b0};
	else if(a[21]) b[51:0] = {a[21:0],30'b0};
	else if(a[20]) b[51:0] = {a[20:0],31'b0};
	
	else if(a[19]) b[51:0] = {a[19:0],32'b0};
	else if(a[18]) b[51:0] = {a[18:0],33'b0};
	else if(a[17]) b[51:0] = {a[17:0],34'b0};
	else if(a[16]) b[51:0] = {a[16:0],35'b0};
	else if(a[15]) b[51:0] = {a[15:0],36'b0};
	else if(a[14]) b[51:0] = {a[14:0],37'b0};
	else if(a[13]) b[51:0] = {a[13:0],38'b0};
	else if(a[12]) b[51:0] = {a[12:0],39'b0};
	else if(a[11]) b[51:0] = {a[11:0],40'b0};
	else if(a[10]) b[51:0] = {a[10:0],41'b0};

	else if(a[9])  b[51:0] = {a[9:0],42'b0};
	else if(a[8])  b[51:0] = {a[8:0],43'b0};
	else if(a[7])  b[51:0] = {a[7:0],44'b0};
	else if(a[6])  b[51:0] = {a[6:0],45'b0};
	else if(a[5])  b[51:0] = {a[5:0],46'b0};
	else if(a[4])  b[51:0] = {a[4:0],47'b0};
	else if(a[3])  b[51:0] = {a[3:0],48'b0};
	else if(a[2])  b[51:0] = {a[2:0],49'b0};
	else if(a[1])  b[51:0] = {a[1:0],50'b0};
	else if(a[0])  b[51:0] = {a[0],51'b0};
	
	else 
		begin
		setzero = 1;
		b = 0;
		end
	
end





endmodule

